`timescale 1ns / 1ps

module level0(
  input  wire [31:0]a,
  input  wire [31:0]b,
  output wire [31:0]p_list,
  output wire [31:0]g_list
);

pg pg_0(a[0], b[0], p_list[0], g_list[0]);
pg pg_1(a[1], b[1], p_list[1], g_list[1]);
pg pg_2(a[2], b[2], p_list[2], g_list[2]);
pg pg_3(a[3], b[3], p_list[3], g_list[3]);
pg pg_4(a[4], b[4], p_list[4], g_list[4]);
pg pg_5(a[5], b[5], p_list[5], g_list[5]);
pg pg_6(a[6], b[6], p_list[6], g_list[6]);
pg pg_7(a[7], b[7], p_list[7], g_list[7]);
pg pg_8(a[8], b[8], p_list[8], g_list[8]);
pg pg_9(a[9], b[9], p_list[9], g_list[9]);
pg pg_10(a[10], b[10], p_list[10], g_list[10]);
pg pg_11(a[11], b[11], p_list[11], g_list[11]);
pg pg_12(a[12], b[12], p_list[12], g_list[12]);
pg pg_13(a[13], b[13], p_list[13], g_list[13]);
pg pg_14(a[14], b[14], p_list[14], g_list[14]);
pg pg_15(a[15], b[15], p_list[15], g_list[15]);
pg pg_16(a[16], b[16], p_list[16], g_list[16]);
pg pg_17(a[17], b[17], p_list[17], g_list[17]);
pg pg_18(a[18], b[18], p_list[18], g_list[18]);
pg pg_19(a[19], b[19], p_list[19], g_list[19]);
pg pg_20(a[20], b[20], p_list[20], g_list[20]);
pg pg_21(a[21], b[21], p_list[21], g_list[21]);
pg pg_22(a[22], b[22], p_list[22], g_list[22]);
pg pg_23(a[23], b[23], p_list[23], g_list[23]);
pg pg_24(a[24], b[24], p_list[24], g_list[24]);
pg pg_25(a[25], b[25], p_list[25], g_list[25]);
pg pg_26(a[26], b[26], p_list[26], g_list[26]);
pg pg_27(a[27], b[27], p_list[27], g_list[27]);
pg pg_28(a[28], b[28], p_list[28], g_list[28]);
pg pg_29(a[29], b[29], p_list[29], g_list[29]);
pg pg_30(a[30], b[30], p_list[30], g_list[30]);
pg pg_31(a[31], b[31], p_list[31], g_list[31]);

endmodule

